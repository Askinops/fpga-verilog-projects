`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.03.2025 04:28:55
// Design Name: 
// Module Name: rotate_right_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rotate_right_32(
    input wire [31:0] a,
    input wire [4:0] amt,
    output reg [31:0] y
    );
    
    
    always @* begin 
        case (amt)
        
        5'd0: y = a;
        5'd1: y = {a[0], a[31:1]};
        5'd2: y = {a[1:0], a[31:2]};
        5'd3: y = {a[2:0], a[31:3]};
        5'd4: y = {a[3:0], a[31:4]};
        5'd5: y = {a[4:0], a[31:5]};
        5'd6: y = {a[5:0], a[31:6]};
        5'd7: y = {a[6:0], a[31:7]};
        5'd8: y = {a[7:0], a[31:8]};
        5'd9: y = {a[8:0], a[31:9]};
        5'd10: y = {a[9:0], a[31:10]};
        5'd11: y = {a[10:0], a[31:11]};
        5'd12: y = {a[11:0], a[31:12]};
        5'd13: y = {a[12:0], a[31:13]};
        5'd14: y = {a[13:0], a[31:14]};
        5'd15: y = {a[14:0], a[31:15]};
        5'd16: y = {a[15:0], a[31:16]};
        5'd17: y = {a[16:0], a[31:17]};
        5'd18: y = {a[17:0], a[31:18]};
        5'd19: y = {a[18:0], a[31:19]};
        5'd20: y = {a[19:0], a[31:20]};
        5'd21: y = {a[20:0], a[31:21]};
        5'd22: y = {a[21:0], a[31:22]};
        5'd23: y = {a[22:0], a[31:23]};
        5'd24: y = {a[23:0], a[31:24]};
        5'd25: y = {a[24:0], a[31:25]};
        5'd26: y = {a[25:0], a[31:26]};
        5'd27: y = {a[26:0], a[31:27]};
        5'd28: y = {a[27:0], a[31:28]};
        5'd29: y = {a[28:0], a[31:29]};
        5'd30: y = {a[29:0], a[31:30]};
        5'd31: y = {a[30:0], a[31]};
        default: y = a;
        
        endcase
    
    
    end 
    
endmodule
